// fir.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module fir (
		input  wire        begin_load_reset_n,   // begin_load.reset_n
		input  wire        clk_clk,              //        clk.clk
		input  wire [18:0] input_data,           //      input.data
		input  wire        input_valid,          //           .valid
		input  wire [1:0]  input_error,          //           .error
		input  wire        input_startofpacket,  //           .startofpacket
		input  wire        input_endofpacket,    //           .endofpacket
		output wire [31:0] output_data,          //     output.data
		output wire        output_valid,         //           .valid
		output wire [1:0]  output_error,         //           .error
		output wire        output_startofpacket, //           .startofpacket
		output wire        output_endofpacket,   //           .endofpacket
		output wire [2:0]  output_channel,       //           .channel
		input  wire        reset_reset_n,        //      reset.reset_n
		input  wire [9:0]  slave_address,        //      slave.address
		input  wire [0:0]  slave_write,          //           .write
		input  wire [15:0] slave_writedata       //           .writedata
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> fir_compiler_ii_0:reset_n

	fir_fir_compiler_ii_0 fir_compiler_ii_0 (
		.clk                (clk_clk),                         //                     clk.clk
		.reset_n            (~rst_controller_reset_out_reset), //                     rst.reset_n
		.ast_sink_data      (input_data),                      //   avalon_streaming_sink.data
		.ast_sink_valid     (input_valid),                     //                        .valid
		.ast_sink_error     (input_error),                     //                        .error
		.ast_sink_sop       (input_startofpacket),             //                        .startofpacket
		.ast_sink_eop       (input_endofpacket),               //                        .endofpacket
		.ast_source_data    (output_data),                     // avalon_streaming_source.data
		.ast_source_valid   (output_valid),                    //                        .valid
		.ast_source_error   (output_error),                    //                        .error
		.ast_source_sop     (output_startofpacket),            //                        .startofpacket
		.ast_source_eop     (output_endofpacket),              //                        .endofpacket
		.ast_source_channel (output_channel),                  //                        .channel
		.coeff_in_clk       (clk_clk),                         //             coeff_clock.clk
		.coeff_in_areset    (begin_load_reset_n),              //             coeff_reset.reset_n
		.coeff_in_address   (slave_address),                   //         avalon_mm_slave.address
		.coeff_in_we        (slave_write),                     //                        .write
		.coeff_in_data      (slave_writedata)                  //                        .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
